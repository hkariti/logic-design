library ieee;
use IEEE.std_logic_1164.all;

entity ContComp is
port (CLK : in std_logic; --Clock, active high
      RSTn : in std_logic --Async. Reset, active low
  );
end entity;

architecture behavior of ContComp is

begin

-- add your code here

end behavior;
